** sch_path: /home/designer/shared/OS_AnalogIC_UCU_July2025/Python_layout/transmission_gate/tgate_inv.sch
.subckt tgate_inv B SEL A VDD_D VSS_D
*.PININFO B:B SEL:B A:B VDD_D:B VSS_D:B
M1 B SEL A VSS_D sg13_lv_nmos l=1u w=0.4u ng=1 m=1
M2 A NSEL B B sg13_lv_pmos l=1u w=1.2u ng=1 m=1
x1 SEL VDD_D VSS_D NSEL sg13g2_inv_1
**** begin user architecture code


*.include '/opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice'

.subckt sg13g2_inv_1 A VDD VSS Y
M1 Y A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M0 Y A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends

**** end user architecture code
.ends
.end
