* Extracted by KLayout with SG13G2 LVS runset on : 02/07/2025 14:23

.SUBCKT tgate_inv
M$1 \$1 \$5 \$4 \$1 sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p PS=2.18u
+ PD=2.18u
M$2 \$6 \$5 \$3 \$1 sg13_lv_nmos L=1u W=0.4u AS=0.136p AD=0.136p PS=1.48u
+ PD=1.48u
M$3 \$2 \$5 \$4 \$2 sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p PS=2.94u
+ PD=2.94u
M$4 \$6 \$4 \$3 \$3 sg13_lv_pmos L=1u W=1.2u AS=0.408p AD=0.408p PS=3.08u
+ PD=3.08u
.ENDS tgate_inv
