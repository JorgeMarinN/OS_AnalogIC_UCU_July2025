** sch_path: /home/designer/shared/OS_AnalogIC_UCU_July2025/Day2/tb_transmission_gate.sch
**.subckt tb_transmission_gate vin1 vout vdd
*.iopin vin1
*.iopin vout
*.iopin vdd
x1 vout GND vdd vin1 vdd GND transmission_gate
x2 vout vdd GND net2 vdd GND transmission_gate
E1 net1 GND vin1 GND 1
vin2 net2 net1 0
**** begin user architecture code


*.param v_max = 1.2
vin1 vin1 0 dc=0.6
vout vout 0 dc=0
vdd vdd 0 dc=1.2

.control
save all

dc vin1 0 1 0.01

meas dc IMAX FIND i(vin2) WHEN vin1=1

plot i(vin1)
plot i(vin2)
let RON = -1/IMAX
print RON


.endc




.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends

* expanding   symbol:  transmission_gate.sym # of pins=6
** sym_path: /home/designer/shared/OS_AnalogIC_UCU_July2025/Day2/transmission_gate.sym
** sch_path: /home/designer/shared/OS_AnalogIC_UCU_July2025/Day2/transmission_gate.sch
.subckt transmission_gate B GN GP A BP BN
*.iopin B
*.iopin GN
*.iopin A
*.iopin GP
*.iopin BN
*.iopin BP
XM1 A GN B BN sg13_lv_nmos w=0.4u l=0.13u ng=1 m=10
XM2 A GP B BP sg13_lv_pmos w=1.2u l=0.13u ng=1 m=10
.ends

.GLOBAL GND
.end
