** sch_path: /home/designer/shared/OS_AnalogIC_UCU_July2025/Day1/tb_inv_1_manual.sch
**.subckt tb_inv_1_manual vin vout vdd
*.iopin vin
*.iopin vout
*.iopin vdd
x1 vdd vin vout GND inv_1_manual
**** begin user architecture code



vin vin 0 dc=0.6
vdd vdd 0 dc=1.2

.control
save all

dc vin 0 1.2 0.01

plot v(vout)


.endc




.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends

* expanding   symbol:  inv_1_manual.sym # of pins=4
** sym_path: /home/designer/shared/OS_AnalogIC_UCU_July2025/Day1/inv_1_manual.sym
** sch_path: /home/designer/shared/OS_AnalogIC_UCU_July2025/Day1/inv_1_manual.sch
.subckt inv_1_manual VDD_D A Y VSS_D
*.iopin VDD_D
*.iopin VSS_D
*.iopin A
*.iopin Y
XM1 VSS_D A Y VSS_D sg13_lv_nmos w=0.74u l=0.13u ng=1 m=1
XM2 Y A VDD_D VDD_D sg13_lv_pmos w=1.12u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
